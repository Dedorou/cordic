module atan_table (
input  logic [ 4 : 0] addr,

output logic [31 : 0] data_o
);

logic [31 : 0] atan_table [0 : 30];
assign atan_table[00] = 'b00100000000000000000000000000000; // 0x20000000 | 45.0000 -> atan(2^0)
assign atan_table[01] = 'b00010010111001000000010100011101; // 0x12e4051d | 26.5651 -> atan(2^-1)
assign atan_table[02] = 'b00001001111110110011100001011011; // 0x09fb385b | 14.0362 -> atan(2^-2)
assign atan_table[03] = 'b00000101000100010001000111010100; // 0x051111d4 |  7.1250 -> atan(2^-3)
assign atan_table[04] = 'b00000010100010110000110101000011; // 0x028b0d43 |  3.5763 -> atan(2^-4)
assign atan_table[05] = 'b00000001010001011101011111100001; // 0x0145d7e1 |  1.7899 -> atan(2^-5)
assign atan_table[06] = 'b00000000101000101111011000011110; // 0x00a2f61e |  0.8952 -> atan(2^-6)
assign atan_table[07] = 'b00000000010100010111110001010101; // 0x00517c55 |  0.4476 -> atan(2^-7)
assign atan_table[08] = 'b00000000001010001011111001010011; // 0x0028be53 |  0.2238 -> atan(2^-8)
assign atan_table[09] = 'b00000000000101000101111100101110; // 0x00145f2e |  0.1119 -> atan(2^-9)
assign atan_table[10] = 'b00000000000010100010111110011000; // 0x000a2f98 |  0.0560 -> atan(2^-10)
assign atan_table[11] = 'b00000000000001010001011111001100; // 0x000517cc |  0.0280 -> atan(2^-11)
assign atan_table[12] = 'b00000000000000101000101111100110; // 0x00028be6 |  0.0140 -> atan(2^-12)
assign atan_table[13] = 'b00000000000000010100010111110011; // 0x000145f3 |  0.0070 -> atan(2^-13)
assign atan_table[14] = 'b00000000000000001010001011111001; // 0x0000a2f9 |  0.0035 -> atan(2^-14)
assign atan_table[15] = 'b00000000000000000101000101111100; // 0x0000517c |  0.0017 -> atan(2^-15)
assign atan_table[16] = 'b00000000000000000010100010111110; // 0x000028be |  0.0009 -> atan(2^-16)
assign atan_table[17] = 'b00000000000000000001010001011111; // 0x0000145f |  0.0004 -> atan(2^-17)
assign atan_table[18] = 'b00000000000000000000101000101111; // 0x00000a2f |  0.0002 -> atan(2^-18)
assign atan_table[19] = 'b00000000000000000000010100010111; // 0x00000517 |  0.0001 -> atan(2^-19)
assign atan_table[20] = 'b00000000000000000000001010001011; // 0x0000028b |  0.0001 -> atan(2^-20)
assign atan_table[21] = 'b00000000000000000000000101000101; // 0x00000145 |  0.0000 -> atan(2^-21)
assign atan_table[22] = 'b00000000000000000000000010100010; // 0x000000a2 |  0.0000 -> atan(2^-22)
assign atan_table[23] = 'b00000000000000000000000001010001; // 0x00000051 |  0.0000 -> atan(2^-23)
assign atan_table[24] = 'b00000000000000000000000000101000; // 0x00000028 |  0.0000 -> atan(2^-24)
assign atan_table[25] = 'b00000000000000000000000000010100; // 0x00000014 |  0.0000 -> atan(2^-25)
assign atan_table[26] = 'b00000000000000000000000000001010; // 0x0000000a |  0.0000 -> atan(2^-26)
assign atan_table[27] = 'b00000000000000000000000000000101; // 0x00000005 |  0.0000 -> atan(2^-27)
assign atan_table[28] = 'b00000000000000000000000000000010; // 0x00000002 |  0.0000 -> atan(2^-28)
assign atan_table[29] = 'b00000000000000000000000000000001; // 0x00000001 |  0.0000 -> atan(2^-29)
assign atan_table[30] = 'b00000000000000000000000000000000; // 0x00000000 |  0.0000 -> atan(2^-30)

assign data_o = atan_table[addr];

endmodule